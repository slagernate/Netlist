; Written by XyceNetlister
; 

; Source File: /home/nates/github/Netlist/examples/spectre_to_xyce/subckts/in.scs
.SUBCKT sub1 d g s b
+ PARAMS: w=60u p1=1000 p2=0.1 vth=0.7 p3={-0.5} p4=1.8 p5=0.7 p6=0.1 p7={-0.02} 

r1 
+ d 
+ g 
+ r=1k 
inst1 
+ d 
+ d1 
+ r={abs(1/w*p1/(1+p2*(v(g,s)-vth-p3*v(b,s)))*(1+pwr(abs(v(d,s)+p6-min(v(d1,s),60))/p4*(1+p7*v(b,s)),p5)))} tc1=0 tc2=0 

.model m1 nmos
+ lmin=0.1u
+ lmax=1.0u
+ wmin=0.5u
+ wmax=10u

.ENDS

