.param vdd = 1.8
.param vss = 0.0
.param width = 1.0u
.param length = 0.18u
.param tox = 4.0n
* Minimal example: Parameter declarations

